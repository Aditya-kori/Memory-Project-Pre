typedef uvm_sequencer#(mem_tx) mem_sequencer;
